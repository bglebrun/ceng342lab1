--------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:   11:19:24 04/10/2018
-- Design Name:
-- Module Name:   C:/Users/7131322/ceng342labs/Lab5/clock_test.vhd
-- Project Name:  Lab5
-- Target Device:
-- Tool versions:
-- Description:
--
-- VHDL Test Bench Created by ISE for module: one_second_clock
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes:
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

ENTITY clock_test IS
END clock_test;

ARCHITECTURE behavior OF clock_test IS

    -- Component Declaration for the Unit Under Test (UUT)

    COMPONENT one_second_clock
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         s_tick : OUT  std_logic
        );
    END COMPONENT;


   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';

 	--Outputs
   signal s_tick : std_logic;

   -- Clock period definitions
   constant clk_period : time := 20 ns;

BEGIN

	-- Instantiate the Unit Under Test (UUT)
   uut: one_second_clock PORT MAP (
          clk => clk,
          reset => reset,
          s_tick => s_tick
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;


   -- Stimulus process
   stim_proc: process
   begin
      -- hold reset state for 100 ns.
      wait for 100 ns;

      wait for clk_period*10;

      -- insert stimulus here

      wait;
   end process;

END;
